library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity GLPLUT2 is 
port(
	inval : in std_logic_vector(7 downto 0);
	outval : out std_logic_vector(7 downto 0)
);

end GLPLUT2;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity GLPLUT3 is 
port(
	inval : in std_logic_vector(7 downto 0);
	outval : out std_logic_vector(7 downto 0)
);

end GLPLUT3;




ARCHITECTURE default of GLPLUT2 is

BEGIN
	 outval<=x"00" when(inval=x"00") else
				x"02" when(inval=x"01") else
				x"04" when(inval=x"02") else
				x"06" when(inval=x"03") else
				x"08" when(inval=x"04") else
				x"0a" when(inval=x"05") else
				x"0c" when(inval=x"06") else
				x"0e" when(inval=x"07") else
				x"10" when(inval=x"08") else
				x"12" when(inval=x"09") else
				x"14" when(inval=x"0a") else
				x"16" when(inval=x"0b") else
				x"18" when(inval=x"0c") else
				x"1a" when(inval=x"0d") else
				x"1c" when(inval=x"0e") else
				x"1e" when(inval=x"0f") else
				x"20" when(inval=x"10") else
				x"22" when(inval=x"11") else
				x"24" when(inval=x"12") else
				x"26" when(inval=x"13") else
				x"28" when(inval=x"14") else
				x"2a" when(inval=x"15") else
				x"2c" when(inval=x"16") else
				x"2e" when(inval=x"17") else
				x"30" when(inval=x"18") else
				x"32" when(inval=x"19") else
				x"34" when(inval=x"1a") else
				x"36" when(inval=x"1b") else
				x"38" when(inval=x"1c") else
				x"3a" when(inval=x"1d") else
				x"3c" when(inval=x"1e") else
				x"3e" when(inval=x"1f") else
				x"40" when(inval=x"20") else
				x"42" when(inval=x"21") else
				x"44" when(inval=x"22") else
				x"46" when(inval=x"23") else
				x"48" when(inval=x"24") else
				x"4a" when(inval=x"25") else
				x"4c" when(inval=x"26") else
				x"4e" when(inval=x"27") else
				x"50" when(inval=x"28") else
				x"52" when(inval=x"29") else
				x"54" when(inval=x"2a") else
				x"56" when(inval=x"2b") else
				x"58" when(inval=x"2c") else
				x"5a" when(inval=x"2d") else
				x"5c" when(inval=x"2e") else
				x"5e" when(inval=x"2f") else
				x"60" when(inval=x"30") else
				x"62" when(inval=x"31") else
				x"64" when(inval=x"32") else
				x"66" when(inval=x"33") else
				x"68" when(inval=x"34") else
				x"6a" when(inval=x"35") else
				x"6c" when(inval=x"36") else
				x"6e" when(inval=x"37") else
				x"70" when(inval=x"38") else
				x"72" when(inval=x"39") else
				x"74" when(inval=x"3a") else
				x"76" when(inval=x"3b") else
				x"78" when(inval=x"3c") else
				x"7a" when(inval=x"3d") else
				x"7c" when(inval=x"3e") else
				x"7e" when(inval=x"3f") else
				x"80" when(inval=x"40") else
				x"82" when(inval=x"41") else
				x"84" when(inval=x"42") else
				x"86" when(inval=x"43") else
				x"88" when(inval=x"44") else
				x"8a" when(inval=x"45") else
				x"8c" when(inval=x"46") else
				x"8e" when(inval=x"47") else
				x"90" when(inval=x"48") else
				x"92" when(inval=x"49") else
				x"94" when(inval=x"4a") else
				x"96" when(inval=x"4b") else
				x"98" when(inval=x"4c") else
				x"9a" when(inval=x"4d") else
				x"9c" when(inval=x"4e") else
				x"9e" when(inval=x"4f") else
				x"a0" when(inval=x"50") else
				x"a2" when(inval=x"51") else
				x"a4" when(inval=x"52") else
				x"a6" when(inval=x"53") else
				x"a8" when(inval=x"54") else
				x"aa" when(inval=x"55") else
				x"ac" when(inval=x"56") else
				x"ae" when(inval=x"57") else
				x"b0" when(inval=x"58") else
				x"b2" when(inval=x"59") else
				x"b4" when(inval=x"5a") else
				x"b6" when(inval=x"5b") else
				x"b8" when(inval=x"5c") else
				x"ba" when(inval=x"5d") else
				x"bc" when(inval=x"5e") else
				x"be" when(inval=x"5f") else
				x"c0" when(inval=x"60") else
				x"c2" when(inval=x"61") else
				x"c4" when(inval=x"62") else
				x"c6" when(inval=x"63") else
				x"c8" when(inval=x"64") else
				x"ca" when(inval=x"65") else
				x"cc" when(inval=x"66") else
				x"ce" when(inval=x"67") else
				x"d0" when(inval=x"68") else
				x"d2" when(inval=x"69") else
				x"d4" when(inval=x"6a") else
				x"d6" when(inval=x"6b") else
				x"d8" when(inval=x"6c") else
				x"da" when(inval=x"6d") else
				x"dc" when(inval=x"6e") else
				x"de" when(inval=x"6f") else
				x"e0" when(inval=x"70") else
				x"e2" when(inval=x"71") else
				x"e4" when(inval=x"72") else
				x"e6" when(inval=x"73") else
				x"e8" when(inval=x"74") else
				x"ea" when(inval=x"75") else
				x"ec" when(inval=x"76") else
				x"ee" when(inval=x"77") else
				x"f0" when(inval=x"78") else
				x"f2" when(inval=x"79") else
				x"f4" when(inval=x"7a") else
				x"f6" when(inval=x"7b") else
				x"f8" when(inval=x"7c") else
				x"fa" when(inval=x"7d") else
				x"fc" when(inval=x"7e") else
				x"fe" when(inval=x"7f") else
				x"1b" when(inval=x"80") else
				x"19" when(inval=x"81") else
				x"1f" when(inval=x"82") else
				x"1d" when(inval=x"83") else
				x"13" when(inval=x"84") else
				x"11" when(inval=x"85") else
				x"17" when(inval=x"86") else
				x"15" when(inval=x"87") else
				x"0b" when(inval=x"88") else
				x"09" when(inval=x"89") else
				x"0f" when(inval=x"8a") else
				x"0d" when(inval=x"8b") else
				x"03" when(inval=x"8c") else
				x"01" when(inval=x"8d") else
				x"07" when(inval=x"8e") else
				x"05" when(inval=x"8f") else
				x"3b" when(inval=x"90") else
				x"39" when(inval=x"91") else
				x"3f" when(inval=x"92") else
				x"3d" when(inval=x"93") else
				x"33" when(inval=x"94") else
				x"31" when(inval=x"95") else
				x"37" when(inval=x"96") else
				x"35" when(inval=x"97") else
				x"2b" when(inval=x"98") else
				x"29" when(inval=x"99") else
				x"2f" when(inval=x"9a") else
				x"2d" when(inval=x"9b") else
				x"23" when(inval=x"9c") else
				x"21" when(inval=x"9d") else
				x"27" when(inval=x"9e") else
				x"25" when(inval=x"9f") else
				x"5b" when(inval=x"a0") else
				x"59" when(inval=x"a1") else
				x"5f" when(inval=x"a2") else
				x"5d" when(inval=x"a3") else
				x"53" when(inval=x"a4") else
				x"51" when(inval=x"a5") else
				x"57" when(inval=x"a6") else
				x"55" when(inval=x"a7") else
				x"4b" when(inval=x"a8") else
				x"49" when(inval=x"a9") else
				x"4f" when(inval=x"aa") else
				x"4d" when(inval=x"ab") else
				x"43" when(inval=x"ac") else
				x"41" when(inval=x"ad") else
				x"47" when(inval=x"ae") else
				x"45" when(inval=x"af") else
				x"7b" when(inval=x"b0") else
				x"79" when(inval=x"b1") else
				x"7f" when(inval=x"b2") else
				x"7d" when(inval=x"b3") else
				x"73" when(inval=x"b4") else
				x"71" when(inval=x"b5") else
				x"77" when(inval=x"b6") else
				x"75" when(inval=x"b7") else
				x"6b" when(inval=x"b8") else
				x"69" when(inval=x"b9") else
				x"6f" when(inval=x"ba") else
				x"6d" when(inval=x"bb") else
				x"63" when(inval=x"bc") else
				x"61" when(inval=x"bd") else
				x"67" when(inval=x"be") else
				x"65" when(inval=x"bf") else
				x"9b" when(inval=x"c0") else
				x"99" when(inval=x"c1") else
				x"9f" when(inval=x"c2") else
				x"9d" when(inval=x"c3") else
				x"93" when(inval=x"c4") else
				x"91" when(inval=x"c5") else
				x"97" when(inval=x"c6") else
				x"95" when(inval=x"c7") else
				x"8b" when(inval=x"c8") else
				x"89" when(inval=x"c9") else
				x"8f" when(inval=x"ca") else
				x"8d" when(inval=x"cb") else
				x"83" when(inval=x"cc") else
				x"81" when(inval=x"cd") else
				x"87" when(inval=x"ce") else
				x"85" when(inval=x"cf") else
				x"bb" when(inval=x"d0") else
				x"b9" when(inval=x"d1") else
				x"bf" when(inval=x"d2") else
				x"bd" when(inval=x"d3") else
				x"b3" when(inval=x"d4") else
				x"b1" when(inval=x"d5") else
				x"b7" when(inval=x"d6") else
				x"b5" when(inval=x"d7") else
				x"ab" when(inval=x"d8") else
				x"a9" when(inval=x"d9") else
				x"af" when(inval=x"da") else
				x"ad" when(inval=x"db") else
				x"a3" when(inval=x"dc") else
				x"a1" when(inval=x"dd") else
				x"a7" when(inval=x"de") else
				x"a5" when(inval=x"df") else
				x"db" when(inval=x"e0") else
				x"d9" when(inval=x"e1") else
				x"df" when(inval=x"e2") else
				x"dd" when(inval=x"e3") else
				x"d3" when(inval=x"e4") else
				x"d1" when(inval=x"e5") else
				x"d7" when(inval=x"e6") else
				x"d5" when(inval=x"e7") else
				x"cb" when(inval=x"e8") else
				x"c9" when(inval=x"e9") else
				x"cf" when(inval=x"ea") else
				x"cd" when(inval=x"eb") else
				x"c3" when(inval=x"ec") else
				x"c1" when(inval=x"ed") else
				x"c7" when(inval=x"ee") else
				x"c5" when(inval=x"ef") else
				x"fb" when(inval=x"f0") else
				x"f9" when(inval=x"f1") else
				x"ff" when(inval=x"f2") else
				x"fd" when(inval=x"f3") else
				x"f3" when(inval=x"f4") else
				x"f1" when(inval=x"f5") else
				x"f7" when(inval=x"f6") else
				x"f5" when(inval=x"f7") else
				x"eb" when(inval=x"f8") else
				x"e9" when(inval=x"f9") else
				x"ef" when(inval=x"fa") else
				x"ed" when(inval=x"fb") else
				x"e3" when(inval=x"fc") else
				x"e1" when(inval=x"fd") else
				x"e7" when(inval=x"fe") else
				x"e5";
END default;



ARCHITECTURE default of GLPLUT3 is

BEGIN
	
	 outval<=x"00" when(inval=x"00") else
				x"03" when(inval=x"01") else
				x"06" when(inval=x"02") else
				x"05" when(inval=x"03") else
				x"0c" when(inval=x"04") else
				x"0f" when(inval=x"05") else
				x"0a" when(inval=x"06") else
				x"09" when(inval=x"07") else
				x"18" when(inval=x"08") else
				x"1b" when(inval=x"09") else
				x"1e" when(inval=x"0a") else
				x"1d" when(inval=x"0b") else
				x"14" when(inval=x"0c") else
				x"17" when(inval=x"0d") else
				x"12" when(inval=x"0e") else
				x"11" when(inval=x"0f") else
				x"30" when(inval=x"10") else
				x"33" when(inval=x"11") else
				x"36" when(inval=x"12") else
				x"35" when(inval=x"13") else
				x"3c" when(inval=x"14") else
				x"3f" when(inval=x"15") else
				x"3a" when(inval=x"16") else
				x"39" when(inval=x"17") else
				x"28" when(inval=x"18") else
				x"2b" when(inval=x"19") else
				x"2e" when(inval=x"1a") else
				x"2d" when(inval=x"1b") else
				x"24" when(inval=x"1c") else
				x"27" when(inval=x"1d") else
				x"22" when(inval=x"1e") else
				x"21" when(inval=x"1f") else
				x"60" when(inval=x"20") else
				x"63" when(inval=x"21") else
				x"66" when(inval=x"22") else
				x"65" when(inval=x"23") else
				x"6c" when(inval=x"24") else
				x"6f" when(inval=x"25") else
				x"6a" when(inval=x"26") else
				x"69" when(inval=x"27") else
				x"78" when(inval=x"28") else
				x"7b" when(inval=x"29") else
				x"7e" when(inval=x"2a") else
				x"7d" when(inval=x"2b") else
				x"74" when(inval=x"2c") else
				x"77" when(inval=x"2d") else
				x"72" when(inval=x"2e") else
				x"71" when(inval=x"2f") else
				x"50" when(inval=x"30") else
				x"53" when(inval=x"31") else
				x"56" when(inval=x"32") else
				x"55" when(inval=x"33") else
				x"5c" when(inval=x"34") else
				x"5f" when(inval=x"35") else
				x"5a" when(inval=x"36") else
				x"59" when(inval=x"37") else
				x"48" when(inval=x"38") else
				x"4b" when(inval=x"39") else
				x"4e" when(inval=x"3a") else
				x"4d" when(inval=x"3b") else
				x"44" when(inval=x"3c") else
				x"47" when(inval=x"3d") else
				x"42" when(inval=x"3e") else
				x"41" when(inval=x"3f") else
				x"c0" when(inval=x"40") else
				x"c3" when(inval=x"41") else
				x"c6" when(inval=x"42") else
				x"c5" when(inval=x"43") else
				x"cc" when(inval=x"44") else
				x"cf" when(inval=x"45") else
				x"ca" when(inval=x"46") else
				x"c9" when(inval=x"47") else
				x"d8" when(inval=x"48") else
				x"db" when(inval=x"49") else
				x"de" when(inval=x"4a") else
				x"dd" when(inval=x"4b") else
				x"d4" when(inval=x"4c") else
				x"d7" when(inval=x"4d") else
				x"d2" when(inval=x"4e") else
				x"d1" when(inval=x"4f") else
				x"f0" when(inval=x"50") else
				x"f3" when(inval=x"51") else
				x"f6" when(inval=x"52") else
				x"f5" when(inval=x"53") else
				x"fc" when(inval=x"54") else
				x"ff" when(inval=x"55") else
				x"fa" when(inval=x"56") else
				x"f9" when(inval=x"57") else
				x"e8" when(inval=x"58") else
				x"eb" when(inval=x"59") else
				x"ee" when(inval=x"5a") else
				x"ed" when(inval=x"5b") else
				x"e4" when(inval=x"5c") else
				x"e7" when(inval=x"5d") else
				x"e2" when(inval=x"5e") else
				x"e1" when(inval=x"5f") else
				x"a0" when(inval=x"60") else
				x"a3" when(inval=x"61") else
				x"a6" when(inval=x"62") else
				x"a5" when(inval=x"63") else
				x"ac" when(inval=x"64") else
				x"af" when(inval=x"65") else
				x"aa" when(inval=x"66") else
				x"a9" when(inval=x"67") else
				x"b8" when(inval=x"68") else
				x"bb" when(inval=x"69") else
				x"be" when(inval=x"6a") else
				x"bd" when(inval=x"6b") else
				x"b4" when(inval=x"6c") else
				x"b7" when(inval=x"6d") else
				x"b2" when(inval=x"6e") else
				x"b1" when(inval=x"6f") else
				x"90" when(inval=x"70") else
				x"93" when(inval=x"71") else
				x"96" when(inval=x"72") else
				x"95" when(inval=x"73") else
				x"9c" when(inval=x"74") else
				x"9f" when(inval=x"75") else
				x"9a" when(inval=x"76") else
				x"99" when(inval=x"77") else
				x"88" when(inval=x"78") else
				x"8b" when(inval=x"79") else
				x"8e" when(inval=x"7a") else
				x"8d" when(inval=x"7b") else
				x"84" when(inval=x"7c") else
				x"87" when(inval=x"7d") else
				x"82" when(inval=x"7e") else
				x"81" when(inval=x"7f") else
				x"9b" when(inval=x"80") else
				x"98" when(inval=x"81") else
				x"9d" when(inval=x"82") else
				x"9e" when(inval=x"83") else
				x"97" when(inval=x"84") else
				x"94" when(inval=x"85") else
				x"91" when(inval=x"86") else
				x"92" when(inval=x"87") else
				x"83" when(inval=x"88") else
				x"80" when(inval=x"89") else
				x"85" when(inval=x"8a") else
				x"86" when(inval=x"8b") else
				x"8f" when(inval=x"8c") else
				x"8c" when(inval=x"8d") else
				x"89" when(inval=x"8e") else
				x"8a" when(inval=x"8f") else
				x"ab" when(inval=x"90") else
				x"a8" when(inval=x"91") else
				x"ad" when(inval=x"92") else
				x"ae" when(inval=x"93") else
				x"a7" when(inval=x"94") else
				x"a4" when(inval=x"95") else
				x"a1" when(inval=x"96") else
				x"a2" when(inval=x"97") else
				x"b3" when(inval=x"98") else
				x"b0" when(inval=x"99") else
				x"b5" when(inval=x"9a") else
				x"b6" when(inval=x"9b") else
				x"bf" when(inval=x"9c") else
				x"bc" when(inval=x"9d") else
				x"b9" when(inval=x"9e") else
				x"ba" when(inval=x"9f") else
				x"fb" when(inval=x"a0") else
				x"f8" when(inval=x"a1") else
				x"fd" when(inval=x"a2") else
				x"fe" when(inval=x"a3") else
				x"f7" when(inval=x"a4") else
				x"f4" when(inval=x"a5") else
				x"f1" when(inval=x"a6") else
				x"f2" when(inval=x"a7") else
				x"e3" when(inval=x"a8") else
				x"e0" when(inval=x"a9") else
				x"e5" when(inval=x"aa") else
				x"e6" when(inval=x"ab") else
				x"ef" when(inval=x"ac") else
				x"ec" when(inval=x"ad") else
				x"e9" when(inval=x"ae") else
				x"ea" when(inval=x"af") else
				x"cb" when(inval=x"b0") else
				x"c8" when(inval=x"b1") else
				x"cd" when(inval=x"b2") else
				x"ce" when(inval=x"b3") else
				x"c7" when(inval=x"b4") else
				x"c4" when(inval=x"b5") else
				x"c1" when(inval=x"b6") else
				x"c2" when(inval=x"b7") else
				x"d3" when(inval=x"b8") else
				x"d0" when(inval=x"b9") else
				x"d5" when(inval=x"ba") else
				x"d6" when(inval=x"bb") else
				x"df" when(inval=x"bc") else
				x"dc" when(inval=x"bd") else
				x"d9" when(inval=x"be") else
				x"da" when(inval=x"bf") else
				x"5b" when(inval=x"c0") else
				x"58" when(inval=x"c1") else
				x"5d" when(inval=x"c2") else
				x"5e" when(inval=x"c3") else
				x"57" when(inval=x"c4") else
				x"54" when(inval=x"c5") else
				x"51" when(inval=x"c6") else
				x"52" when(inval=x"c7") else
				x"43" when(inval=x"c8") else
				x"40" when(inval=x"c9") else
				x"45" when(inval=x"ca") else
				x"46" when(inval=x"cb") else
				x"4f" when(inval=x"cc") else
				x"4c" when(inval=x"cd") else
				x"49" when(inval=x"ce") else
				x"4a" when(inval=x"cf") else
				x"6b" when(inval=x"d0") else
				x"68" when(inval=x"d1") else
				x"6d" when(inval=x"d2") else
				x"6e" when(inval=x"d3") else
				x"67" when(inval=x"d4") else
				x"64" when(inval=x"d5") else
				x"61" when(inval=x"d6") else
				x"62" when(inval=x"d7") else
				x"73" when(inval=x"d8") else
				x"70" when(inval=x"d9") else
				x"75" when(inval=x"da") else
				x"76" when(inval=x"db") else
				x"7f" when(inval=x"dc") else
				x"7c" when(inval=x"dd") else
				x"79" when(inval=x"de") else
				x"7a" when(inval=x"df") else
				x"3b" when(inval=x"e0") else
				x"38" when(inval=x"e1") else
				x"3d" when(inval=x"e2") else
				x"3e" when(inval=x"e3") else
				x"37" when(inval=x"e4") else
				x"34" when(inval=x"e5") else
				x"31" when(inval=x"e6") else
				x"32" when(inval=x"e7") else
				x"23" when(inval=x"e8") else
				x"20" when(inval=x"e9") else
				x"25" when(inval=x"ea") else
				x"26" when(inval=x"eb") else
				x"2f" when(inval=x"ec") else
				x"2c" when(inval=x"ed") else
				x"29" when(inval=x"ee") else
				x"2a" when(inval=x"ef") else
				x"0b" when(inval=x"f0") else
				x"08" when(inval=x"f1") else
				x"0d" when(inval=x"f2") else
				x"0e" when(inval=x"f3") else
				x"07" when(inval=x"f4") else
				x"04" when(inval=x"f5") else
				x"01" when(inval=x"f6") else
				x"02" when(inval=x"f7") else
				x"13" when(inval=x"f8") else
				x"10" when(inval=x"f9") else
				x"15" when(inval=x"fa") else
				x"16" when(inval=x"fb") else
				x"1f" when(inval=x"fc") else
				x"1c" when(inval=x"fd") else
				x"19" when(inval=x"fe") else
				x"1a";
end default;
