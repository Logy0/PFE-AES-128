-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_bidir 

-- ============================================================
-- File Name: IOBuff.vhd
-- Megafunction Name(s):
-- 			altiobuf_bidir
--
-- Simulation Library Files(s):
-- 			cycloneiii
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altiobuf_bidir CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone III" ENABLE_BUS_HOLD="FALSE" NUMBER_OF_CHANNELS=128 OPEN_DRAIN_OUTPUT="FALSE" USE_DIFFERENTIAL_MODE="FALSE" USE_DYNAMIC_TERMINATION_CONTROL="FALSE" USE_TERMINATION_CONTROL="FALSE" datain dataio dataout oe
--VERSION_BEGIN 13.1 cbx_altiobuf_bidir 2013:10:23:18:05:48:SJ cbx_mgl 2013:10:23:18:06:54:SJ cbx_stratixiii 2013:10:23:18:05:48:SJ cbx_stratixv 2013:10:23:18:05:48:SJ  VERSION_END

 LIBRARY cycloneiii;
 USE cycloneiii.all;

--synthesis_resources = cycloneiii_io_ibuf 128 cycloneiii_io_obuf 128 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  IOBuff_iobuf_bidir_42p IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (127 DOWNTO 0);
		 dataio	:	INOUT  STD_LOGIC_VECTOR (127 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (127 DOWNTO 0);
		 oe	:	IN  STD_LOGIC_VECTOR (127 DOWNTO 0)
	 ); 
 END IOBuff_iobuf_bidir_42p;

 ARCHITECTURE RTL OF IOBuff_iobuf_bidir_42p IS

	 SIGNAL  wire_ibufa_i	:	STD_LOGIC_VECTOR (127 DOWNTO 0);
	 SIGNAL  wire_ibufa_o	:	STD_LOGIC_VECTOR (127 DOWNTO 0);
	 SIGNAL  wire_obufa_i	:	STD_LOGIC_VECTOR (127 DOWNTO 0);
	 SIGNAL  wire_obufa_o	:	STD_LOGIC_VECTOR (127 DOWNTO 0);
	 SIGNAL  wire_obufa_oe	:	STD_LOGIC_VECTOR (127 DOWNTO 0);
	 COMPONENT  cycloneiii_io_ibuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		differential_mode	:	STRING := "false";
		simulate_z_as	:	STRING := "Z";
		lpm_type	:	STRING := "cycloneiii_io_ibuf"
	 );
	 PORT
	 ( 
		i	:	IN STD_LOGIC := '0';
		ibar	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiii_io_obuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		open_drain_output	:	STRING := "false";
		lpm_type	:	STRING := "cycloneiii_io_obuf"
	 );
	 PORT
	 ( 
		i	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC;
		obar	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		seriesterminationcontrol	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	dataio <= wire_obufa_o;
	dataout <= wire_ibufa_o;
	wire_ibufa_i <= dataio;
	loop0 : FOR i IN 0 TO 127 GENERATE 
	  ibufa :  cycloneiii_io_ibuf
	  GENERIC MAP (
		bus_hold => "false",
		differential_mode => "false"
	  )
	  PORT MAP ( 
		i => wire_ibufa_i(i),
		o => wire_ibufa_o(i)
	  );
	END GENERATE loop0;
	wire_obufa_i <= datain;
	wire_obufa_oe <= oe;
	loop1 : FOR i IN 0 TO 127 GENERATE 
	  obufa :  cycloneiii_io_obuf
	  GENERIC MAP (
		bus_hold => "false",
		open_drain_output => "false"
	  )
	  PORT MAP ( 
		i => wire_obufa_i(i),
		o => wire_obufa_o(i),
		oe => wire_obufa_oe(i)
	  );
	END GENERATE loop1;

 END RTL; --IOBuff_iobuf_bidir_42p
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY IOBuff IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		oe		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		dataio		: INOUT STD_LOGIC_VECTOR (127 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (127 DOWNTO 0)
	);
END IOBuff;


ARCHITECTURE RTL OF iobuff IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (127 DOWNTO 0);



	COMPONENT IOBuff_iobuf_bidir_42p
	PORT (
			datain	: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
			dataio	: INOUT STD_LOGIC_VECTOR (127 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (127 DOWNTO 0);
			oe	: IN STD_LOGIC_VECTOR (127 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(127 DOWNTO 0);

	IOBuff_iobuf_bidir_42p_component : IOBuff_iobuf_bidir_42p
	PORT MAP (
		datain => datain,
		oe => oe,
		dataout => sub_wire0,
		dataio => dataio
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "128"
-- Retrieval info: CONSTANT: open_drain_output STRING "FALSE"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_dynamic_termination_control STRING "FALSE"
-- Retrieval info: CONSTANT: use_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 128 0 INPUT NODEFVAL "datain[127..0]"
-- Retrieval info: USED_PORT: dataio 0 0 128 0 BIDIR NODEFVAL "dataio[127..0]"
-- Retrieval info: USED_PORT: dataout 0 0 128 0 OUTPUT NODEFVAL "dataout[127..0]"
-- Retrieval info: USED_PORT: oe 0 0 128 0 INPUT NODEFVAL "oe[127..0]"
-- Retrieval info: CONNECT: @datain 0 0 128 0 datain 0 0 128 0
-- Retrieval info: CONNECT: @oe 0 0 128 0 oe 0 0 128 0
-- Retrieval info: CONNECT: dataio 0 0 128 0 @dataio 0 0 128 0
-- Retrieval info: CONNECT: dataout 0 0 128 0 @dataout 0 0 128 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL IOBuff.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL IOBuff.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL IOBuff.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL IOBuff.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL IOBuff_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cycloneiii
