library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity Sbox is 
port(
		input : in std_logic_vector(7 downto 0);
		out_data : out std_logic_vector(7 downto 0)		
);
end Sbox;


architecture sbox_arch of Sbox is 


begin	
	  --out_data<=input;
	  
	  with input select out_data<=
				   x"63" when x"00",
					x"7c" when x"01",
					x"77" when x"02",
					x"7b" when x"03",
					x"f2" when x"04",
					x"6b" when x"05",
					x"6f" when x"06",
					x"c5" when x"07",
					x"30" when x"08",
					x"01" when x"09",
					x"67" when x"0a",
					x"2b" when x"0b",
					x"fe" when x"0c",
					x"d7" when x"0d",
					x"ab" when x"0e",
					x"76" when x"0f",
					x"ca" when x"10",
					x"82" when x"11",
					x"c9" when x"12",
					x"7d" when x"13",
					x"fa" when x"14",
					x"59" when x"15",
					x"47" when x"16",
					x"f0" when x"17",
					x"ad" when x"18",
					x"d4" when x"19",
					x"a2" when x"1a",
					x"af" when x"1b",
					x"9c" when x"1c",
					x"a4" when x"1d",
					x"72" when x"1e",
					x"c0" when x"1f",
					x"b7" when x"20",
					x"fd" when x"21",
					x"93" when x"22",
					x"26" when x"23",
					x"36" when x"24",
					x"3f" when x"25",
					x"f7" when x"26",
					x"cc" when x"27",
					x"34" when x"28",
					x"a5" when x"29",
					x"e5" when x"2a",
					x"f1" when x"2b",
					x"71" when x"2c",
					x"d8" when x"2d",
					x"31" when x"2e",
					x"15" when x"2f",
					x"04" when x"30",
					x"c7" when x"31",
					x"23" when x"32",
					x"c3" when x"33",
					x"18" when x"34",
					x"96" when x"35",
					x"05" when x"36",
					x"9a" when x"37",
					x"07" when x"38",
					x"12" when x"39",
					x"80" when x"3a",
					x"e2" when x"3b",
					x"eb" when x"3c",
					x"27" when x"3d",
					x"b2" when x"3e",
					x"75" when x"3f",
					x"09" when x"40",
					x"83" when x"41",
					x"2c" when x"42",
					x"1a" when x"43",
					x"1b" when x"44",
					x"6e" when x"45",
					x"5a" when x"46",
					x"a0" when x"47",
					x"52" when x"48",
					x"3b" when x"49",
					x"d6" when x"4a",
					x"b3" when x"4b",
					x"29" when x"4c",
					x"e3" when x"4d",
					x"2f" when x"4e",
					x"84" when x"4f",
					x"53" when x"50",
					x"d1" when x"51",
					x"00" when x"52",
					x"ed" when x"53",
					x"20" when x"54",
					x"fc" when x"55",
					x"b1" when x"56",
					x"5b" when x"57",
					x"6a" when x"58",
					x"cb" when x"59",
					x"be" when x"5a",
					x"39" when x"5b",
					x"4a" when x"5c",
					x"4c" when x"5d",
					x"58" when x"5e",
					x"cf" when x"5f",
					x"d0" when x"60",
					x"ef" when x"61",
					x"aa" when x"62",
					x"fb" when x"63",
					x"43" when x"64",
					x"4d" when x"65",
					x"33" when x"66",
					x"85" when x"67",
					x"45" when x"68",
					x"f9" when x"69",
					x"02" when x"6a",
					x"7f" when x"6b",
					x"50" when x"6c",
					x"3c" when x"6d",
					x"9f" when x"6e",
					x"a8" when x"6f",
					x"51" when x"70",
					x"a3" when x"71",
					x"40" when x"72",
					x"8f" when x"73",
					x"92" when x"74",
					x"9d" when x"75",
					x"38" when x"76",
					x"f5" when x"77",
					x"bc" when x"78",
					x"b6" when x"79",
					x"da" when x"7a",
					x"21" when x"7b",
					x"10" when x"7c",
					x"ff" when x"7d",
					x"f3" when x"7e",
					x"d2" when x"7f",
					x"cd" when x"80",
					x"0c" when x"81",
					x"13" when x"82",
					x"ec" when x"83",
					x"5f" when x"84",
					x"97" when x"85",
					x"44" when x"86",
					x"17" when x"87",
					x"c4" when x"88",
					x"a7" when x"89",
					x"7e" when x"8a",
					x"3d" when x"8b",
					x"64" when x"8c",
					x"5d" when x"8d",
					x"19" when x"8e",
					x"73" when x"8f",
					x"60" when x"90",
					x"81" when x"91",
					x"4f" when x"92",
					x"dc" when x"93",
					x"22" when x"94",
					x"2a" when x"95",
					x"90" when x"96",
					x"88" when x"97",
					x"46" when x"98",
					x"ee" when x"99",
					x"b8" when x"9a",
					x"14" when x"9b",
					x"de" when x"9c",
					x"5e" when x"9d",
					x"0b" when x"9e",
					x"db" when x"9f",
					x"e0" when x"a0",
					x"32" when x"a1",
					x"3a" when x"a2",
					x"0a" when x"a3",
					x"49" when x"a4",
					x"06" when x"a5",
					x"24" when x"a6",
					x"5c" when x"a7",
					x"c2" when x"a8",
					x"d3" when x"a9",
					x"ac" when x"aa",
					x"62" when x"ab",
					x"91" when x"ac",
					x"95" when x"ad",
					x"e4" when x"ae",
					x"79" when x"af",
					x"e7" when x"b0",
					x"c8" when x"b1",
					x"37" when x"b2",
					x"6d" when x"b3",
					x"8d" when x"b4",
					x"d5" when x"b5",
					x"4e" when x"b6",
					x"a9" when x"b7",
					x"6c" when x"b8",
					x"56" when x"b9",
					x"f4" when x"ba",
					x"ea" when x"bb",
					x"65" when x"bc",
					x"7a" when x"bd",
					x"ae" when x"be",
					x"08" when x"bf",
					x"ba" when x"c0",
					x"78" when x"c1",
					x"25" when x"c2",
					x"2e" when x"c3",
					x"1c" when x"c4",
					x"a6" when x"c5",
					x"b4" when x"c6",
					x"c6" when x"c7",
					x"e8" when x"c8",
					x"dd" when x"c9",
					x"74" when x"ca",
					x"1f" when x"cb",
					x"4b" when x"cc",
					x"bd" when x"cd",
					x"8b" when x"ce",
					x"8a" when x"cf",
					x"70" when x"d0",
					x"3e" when x"d1",
					x"b5" when x"d2",
					x"66" when x"d3",
					x"48" when x"d4",
					x"03" when x"d5",
					x"f6" when x"d6",
					x"0e" when x"d7",
					x"61" when x"d8",
					x"35" when x"d9",
					x"57" when x"da",
					x"b9" when x"db",
					x"86" when x"dc",
					x"c1" when x"dd",
					x"1d" when x"de",
					x"9e" when x"df",
					x"e1" when x"e0",
					x"f8" when x"e1",
					x"98" when x"e2",
					x"11" when x"e3",
					x"69" when x"e4",
					x"d9" when x"e5",
					x"8e" when x"e6",
					x"94" when x"e7",
					x"9b" when x"e8",
					x"1e" when x"e9",
					x"87" when x"ea",
					x"e9" when x"eb",
					x"ce" when x"ec",
					x"55" when x"ed",
					x"28" when x"ee",
					x"df" when x"ef",
					x"8c" when x"f0",
					x"a1" when x"f1",
					x"89" when x"f2",
					x"0d" when x"f3",
					x"bf" when x"f4",
					x"e6" when x"f5",
					x"42" when x"f6",
					x"68" when x"f7",
					x"41" when x"f8",
					x"99" when x"f9",
					x"2d" when x"fa",
					x"0f" when x"fb",
					x"b0" when x"fc",
					x"54" when x"fd",
					x"bb" when x"fe",
					x"16" when x"ff";
	
end sbox_arch;
